** Profile: "SCHEMATIC1-CASE2_F_400kHz_SIM"  [ C:\Users\elvis\Documents\CSUN\2021-2022\Fall-2021\ECE442L\Lab 2\CMOS-Two-Input-NAND-Gate-Design\ECE442L_ElvisChino-Islas_Lab_2_Case_2_f_400kHz_Pspice_circuit-PSpiceFiles\SCHEMATIC1\CASE2_F_400kHz_SIM.sim ] 

** Creating circuit file "CASE2_F_400kHz_SIM.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../ece442l_elvischino-islas_lab_2_case_2_f_400khz_pspice_circuit-pspicefiles/ece442l_elvischino-islas_lab_2_case_2_f_40"
+ "0khz_pspice_circuit.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 7.5us 0 1ns 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
